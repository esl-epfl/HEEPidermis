// Copyright 2022 EPFL and Politecnico di Torino.
// Solderpad Hardware License, Version 2.1, see LICENSE.md for details.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// File: vref_pkg.sv
// Author: Juan Sapriza
// Date: 26/04/2025
// Description: Package containing definitions for the vREF.

package vref_pkg;

    parameter int unsigned VrefCalibrationWidth = 5;

endpackage
